library verilog;
use verilog.vl_types.all;
entity toplayicidisplay_vlg_vec_tst is
end toplayicidisplay_vlg_vec_tst;
