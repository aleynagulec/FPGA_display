library verilog;
use verilog.vl_types.all;
entity aaa_vlg_vec_tst is
end aaa_vlg_vec_tst;
