library verilog;
use verilog.vl_types.all;
entity toplayici_vlg_vec_tst is
end toplayici_vlg_vec_tst;
