library verilog;
use verilog.vl_types.all;
entity toplayici_vlg_check_tst is
    port(
        cikis0          : in     vl_logic;
        cikis1          : in     vl_logic;
        cikis2          : in     vl_logic;
        cikis3          : in     vl_logic;
        Cout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end toplayici_vlg_check_tst;
